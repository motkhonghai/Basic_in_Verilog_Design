module logicGateUsingGateLevelModel(input );
	and 
endmodule
