/*
+-----+-----+-----+-------+-------------+
|  A  |  B  | Cin |  S    | C_out       |
+-----+-----+-----+-------+-------------+
|  0  |  0  |  0  |   0   |     0       |
+-----+-----+-----+-------+-------------+
|  0  |  0  |  1  |   1   |     0       |
+-----+-----+-----+-------+-------------+
|  0  |  1  |  0  |   1   |     0       |
+-----+-----+-----+-------+-------------+
|  0  |  1  |  1  |   0   |     1       |
+-----+-----+-----+-------+-------------+
|  1  |  0  |  0  |   1   |     0       |
+-----+-----+-----+-------+-------------+
|  1  |  0  |  1  |   0   |     1       |
+-----+-----+-----+-------+-------------+
|  1  |  1  |  0  |   0   |     1       |
+-----+-----+-----+-------+-------------+
|  1  |  1  |  1  |   1   |     1       |
+-----+-----+-----+-------+-------------+

sum = a^b^c
cout = (a&b) + ((a^b)&c)
*/

module full_adder(input a, b, cin, output sum, cout);
    
    wire s1,c1,c2;

    half_adder ha1(a, b, s1, c1);
    half_adder ha2(s1, cin, sum, c2);

    assign cout = c1|c2;
endmodule