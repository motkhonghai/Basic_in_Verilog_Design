/*
+-----+-----+-----+-------+-------------+
|  A  |  B  | Cin |  S    | C_out       |
+-----+-----+-----+-------+-------------+
|  0  |  0  |  0  |   0   |     0       |
+-----+-----+-----+-------+-------------+
|  0  |  0  |  1  |   1   |     0       |
+-----+-----+-----+-------+-------------+
|  0  |  1  |  0  |   1   |     0       |
+-----+-----+-----+-------+-------------+
|  0  |  1  |  1  |   0   |     1       |
+-----+-----+-----+-------+-------------+
|  1  |  0  |  0  |   1   |     0       |
+-----+-----+-----+-------+-------------+
|  1  |  0  |  1  |   0   |     1       |
+-----+-----+-----+-------+-------------+
|  1  |  1  |  0  |   0   |     1       |
+-----+-----+-----+-------+-------------+
|  1  |  1  |  1  |   1   |     1       |
+-----+-----+-----+-------+-------------+

sum = a^b^c
cout = (a&b) | (a&c) | (b&c)
*/

module full_adder(input a, b, cin, output sum, cout);
	assign sum 	= a^b^cin;
	assign cout	= (a&b) | (a&cin) | (b&cin);
endmodule
